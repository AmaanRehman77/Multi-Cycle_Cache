package tb_mp_cache_pkg;
    import uvm_pkg::*;
    `include "uvm_macros.svh"

    `include "tb_mp_cache_params.svh"
    `include "tb_mp_cache_transaction.svh"
    `include "tb_mp_cache_cfg.svh"
    `include "tb_mp_cache_sqr.svh"
    `include "tb_mp_cache_seq.svh"
    `include "tb_mp_cache_driver.svh"
    `include "tb_mp_cache_monitor.svh"
    `include "tb_mp_cache_agent.svh"
    `include "tb_mp_cache_reference_model.svh"
    `include "tb_mp_cache_env.svh"
    `include "tb_mp_cache_test.svh"
    `include "tb_mp_cache_scoreboard.svh"


endpackage : tb_mp_cache_pkg